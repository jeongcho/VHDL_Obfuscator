LIBRARY IEEE; USE IEEE.std_logic_1164.ALL; USE IEEE.std_logic_unsigned.ALL; USE IEEE.numeric_std.ALL; Library UNISIM; use UNISIM.vcomponents.all; entity ADC12020 is Port ( ff66634b612f4d46776431426239796e69595a575831413d3d : in std_logic; ff5265546f48666357584236504c5951756c496d4859773d3d : in std_logic; ff35486432672f59566a33374f395741557145392b47413d3d : in std_logic; ff44636a2f325a3379446b685a472b78523636656767513d3d : in std_logic_vector(11 downto 0); ff3733516e4872384b2b4d313778654b617332752f32413d3d : in std_logic; ff6e3536516f646f71694a6d4152536d735a78574475773d3d : in std_logic_vector(5 downto 0); ff507a534d467a36562f345a534e5755745574326668773d3d : in std_logic_vector(1 downto 0); ff734375372b7345675871315954415046687a5046356b45354d79796e5a506d70346e7835483537776a52733d : in std_logic_vector(1 downto 0); ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d : in std_logic; ff35345579546249415444475676365976357270794f706466634b6948397a6f7466675938636851536461593d : in std_logic; ff35345579546249415444475676365976357270794f754e5335735975446a484354684b506d6d344f6554453d : in std_logic; ff78367278306164782f62776f386552346a615a594c673d3d : out std_logic; ff4f4e713355624a533343352b346e33756246377338673d3d : out std_logic; ff526a78674d6b6743434d707672794536766e71794c513d3d : in std_logic; ff547151597569774e3243584579796a57764a7a6c39673d3d : out std_logic; ff3749554e2f736346657730416b38716a732b745371513d3d : out std_logic; ff545336484f3169516e614c77456c316d622f53482f673d3d : out std_logic; ff336c46794e7a665a41773233795930316930313174513d3d : out std_logic_vector(15 downto 0) ); end ADC12020; architecture Behavioral of ADC12020 is attribute IOB : string; type ff4463694d6d3674306b327471514e62734244666268773d3d is (st_idle, st_line_ave0, st_line_ave1, st_line_ave2, st_line_ave3, st_line_ave4, st_wr0, st_wr1, st_done); signal ff3332356d7477754d64456339442f2b5a6c44727579413d3d : ff4463694d6d3674306b327471514e62734244666268773d3d := st_idle; signal ff6d79702b36614f2b55594a797369344e6c56482b65413d3d : STD_LOGIC_VECTOR(11 downto 0) := (others => '0'); attribute IOB of ff6d79702b36614f2b55594a797369344e6c56482b65413d3d : signal is "TRUE"; signal ff70553469356248674669474e4f396e764b594b7958773d3d : std_logic := '0'; signal ff764d71614b5443474d507a536f41756f6a356a5638773d3d : std_logic := '0'; signal ff6f6f49524b56444d77713077545a545663315a5045413d3d : std_logic_vector(5 downto 0) := (others => '0'); signal ff566578526b744538644b49392b59753658356a6359413d3d : std_logic_vector(7 downto 0) := (others => '0'); signal ff556c7542746b515351533838686b37614254365847513d3d : std_logic := '0'; signal ff5343306145363166474e5241315a39645a6a6d4879773d3d : std_logic := '0'; signal ff71444670796c6e74686577476451676d39424a302f513d3d : std_logic_vector(16 downto 0) := (others => '0'); signal ff49596952527246685a316551654f564e6635662f39413d3d : std_logic_vector(16 downto 0); signal ff74434b38614a354247676547696a3048776554796f513d3d : std_logic := '0'; signal ff4a644751576c526f685a63496b69594a7172304848673d3d : std_logic := '0'; signal ff557746415069796532515158714d554e6632366b38513d3d : std_logic_vector(16 downto 0) := (others => '0'); signal ff644e52654c42493575715935704d6a745041723146773d3d : std_logic_vector(16 downto 0); signal ff463171634a63344666425a514c56473549496f6a35773d3d : std_logic_vector(15 downto 0) := (others => '0'); signal ff366e677746596c337243586a4d5452644a775a4c65673d3d : STD_LOGIC_VECTOR(0 downto 0) := "0"; signal ff6c6475433641737731515947564b576b796a6c6b4c773d3d : STD_LOGIC_VECTOR(13 downto 0) := (others => '0'); signal ff2f4636662f6c3072673535706e41485a3762646854513d3d : std_logic_vector(16 downto 0) := (others => '0'); signal ff714f412b3968364e7561522b464c4e355a4a445231673d3d : std_logic_vector(11 downto 0); signal ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d : std_logic := '0'; signal ff63705a6d713032797a6f6c39647875556a4737556b5545354d79796e5a506d70346e7835483537776a52733d : std_logic := '0'; signal ff41734f64796e456c5746356d69726979457351574d513d3d : STD_LOGIC_VECTOR(13 downto 0); signal ff71696d73453179677739397a633754775874385361773d3d : STD_LOGIC_VECTOR(15 downto 0); signal ff6c52395545616841562b5330335664716b697a3933706466634b6948397a6f7466675938636851536461593d : std_logic; signal ff6c52395545616841562b5330335664716b697a3933754e5335735975446a484354684b506d6d344f6554453d : std_logic; signal ff416f464a616f72316f6c5653574451334b42425836513d3d : std_logic; signal ff364237545642476634566358363657586b6d2b5330673d3d : std_logic_vector(15 downto 0); signal ff442f5a372f344d4f50427876662b55446d74477771673d3d : std_logic := '0'; signal ff64684b35757841614e684d304243786e335a6a5438513d3d : std_logic_vector(15 downto 0) := (others => '0'); signal ff6947484f5a464e57314e6d57485976714235554f44773d3d : std_logic := '0'; signal ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d : std_logic_vector(15 downto 0) := x"A003"; begin process(ff66634b612f4d46776431426239796e69595a575831413d3d) is begin if rising_edge(ff66634b612f4d46776431426239796e69595a575831413d3d) then ff6d79702b36614f2b55594a797369344e6c56482b65413d3d <= ff44636a2f325a3379446b685a472b78523636656767513d3d; end if; end process; process(ff66634b612f4d46776431426239796e69595a575831413d3d) is begin if rising_edge(ff66634b612f4d46776431426239796e69595a575831413d3d) then ff764d71614b5443474d507a536f41756f6a356a5638773d3d <= ff70553469356248674669474e4f396e764b594b7958773d3d; case ff3332356d7477754d64456339442f2b5a6c44727579413d3d is when st_idle => ff70553469356248674669474e4f396e764b594b7958773d3d <= '0'; if (ff3733516e4872384b2b4d313778654b617332752f32413d3d = '1') then if (ff6e3536516f646f71694a6d4152536d735a78574475773d3d /= 0) then if (ff6e3536516f646f71694a6d4152536d735a78574475773d3d - '1' /= ff6f6f49524b56444d77713077545a545663315a5045413d3d) then ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_line_ave0; else ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_line_ave3; end if; else ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_wr0; end if; end if; when st_line_ave0 => ff566578526b744538644b49392b59753658356a6359413d3d <= ff566578526b744538644b49392b59753658356a6359413d3d + '1'; if (ff6f6f49524b56444d77713077545a545663315a5045413d3d = 0) then if (ff566578526b744538644b49392b59753658356a6359413d3d = 1) then ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_line_ave1; ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '0'; ff4a644751576c526f685a63496b69594a7172304848673d3d <= '0'; ff566578526b744538644b49392b59753658356a6359413d3d <= (others => '0'); end if; else if (ff566578526b744538644b49392b59753658356a6359413d3d = 1) then ff566578526b744538644b49392b59753658356a6359413d3d <= (others => '0'); ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_line_ave2; end if; if (ff6f6f49524b56444d77713077545a545663315a5045413d3d(0) = '1') then ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '1'; ff4a644751576c526f685a63496b69594a7172304848673d3d <= '0'; else ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '0'; ff4a644751576c526f685a63496b69594a7172304848673d3d <= '1'; end if; end if; when st_line_ave1 => ff463171634a63344666425a514c56473549496f6a35773d3d <= ff463171634a63344666425a514c56473549496f6a35773d3d + '1'; if (ff463171634a63344666425a514c56473549496f6a35773d3d = 5120) then ff463171634a63344666425a514c56473549496f6a35773d3d <= (others => '0'); ff556c7542746b515351533838686b37614254365847513d3d <= '0'; ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_done; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '1'; else ff556c7542746b515351533838686b37614254365847513d3d <= '1'; ff71444670796c6e74686577476451676d39424a302f513d3d <= "00000" & ff6d79702b36614f2b55594a797369344e6c56482b65413d3d; end if; when st_line_ave2 => ff463171634a63344666425a514c56473549496f6a35773d3d <= ff463171634a63344666425a514c56473549496f6a35773d3d + '1'; ff71444670796c6e74686577476451676d39424a302f513d3d <= ff644e52654c42493575715935704d6a745041723146773d3d + ff6d79702b36614f2b55594a797369344e6c56482b65413d3d; ff557746415069796532515158714d554e6632366b38513d3d <= ff49596952527246685a316551654f564e6635662f39413d3d + ff6d79702b36614f2b55594a797369344e6c56482b65413d3d; if (ff463171634a63344666425a514c56473549496f6a35773d3d = 5198) then ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '0'; ff4a644751576c526f685a63496b69594a7172304848673d3d <= '0'; elsif (ff463171634a63344666425a514c56473549496f6a35773d3d = 5120) then ff463171634a63344666425a514c56473549496f6a35773d3d <= (others => '0'); ff556c7542746b515351533838686b37614254365847513d3d <= '0'; ff74434b38614a354247676547696a3048776554796f513d3d <= '0'; ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '0'; ff4a644751576c526f685a63496b69594a7172304848673d3d <= '0'; ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_done; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '1'; elsif (ff6f6f49524b56444d77713077545a545663315a5045413d3d(0) = '1') then ff556c7542746b515351533838686b37614254365847513d3d <= '0'; ff74434b38614a354247676547696a3048776554796f513d3d <= '1'; elsif (ff6f6f49524b56444d77713077545a545663315a5045413d3d(0) = '0') then ff556c7542746b515351533838686b37614254365847513d3d <= '1'; ff74434b38614a354247676547696a3048776554796f513d3d <= '0'; end if; when st_line_ave3 => ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '1'; ff566578526b744538644b49392b59753658356a6359413d3d <= ff566578526b744538644b49392b59753658356a6359413d3d + '1'; if (ff566578526b744538644b49392b59753658356a6359413d3d = 1) then ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_line_ave4; ff566578526b744538644b49392b59753658356a6359413d3d <= (others => '0'); end if; when st_line_ave4 => ff366e677746596c337243586a4d5452644a775a4c65673d3d <= "1"; ff2f4636662f6c3072673535706e41485a3762646854513d3d <= ff49596952527246685a316551654f564e6635662f39413d3d + ff6d79702b36614f2b55594a797369344e6c56482b65413d3d; if (ff6c6475433641737731515947564b576b796a6c6b4c773d3d = 5117) then ff5343306145363166474e5241315a39645a6a6d4879773d3d <= '0'; ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= ff6c6475433641737731515947564b576b796a6c6b4c773d3d + '1'; elsif (ff6c6475433641737731515947564b576b796a6c6b4c773d3d = 5119) then ff366e677746596c337243586a4d5452644a775a4c65673d3d <= "0"; ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= (others => '0'); ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_done; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '1'; elsif (ff366e677746596c337243586a4d5452644a775a4c65673d3d = "1") then ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= ff6c6475433641737731515947564b576b796a6c6b4c773d3d + '1'; end if; when st_wr0 => ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_wr1; when st_wr1 => ff366e677746596c337243586a4d5452644a775a4c65673d3d <= "1"; if (ff6c6475433641737731515947564b576b796a6c6b4c773d3d = 5119) then ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= (others => '0'); ff366e677746596c337243586a4d5452644a775a4c65673d3d <= "0"; ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_done; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '1'; elsif (ff366e677746596c337243586a4d5452644a775a4c65673d3d = "1") then ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= ff6c6475433641737731515947564b576b796a6c6b4c773d3d + '1'; end if; when st_done => ff556c7542746b515351533838686b37614254365847513d3d <= '0'; ff74434b38614a354247676547696a3048776554796f513d3d <= '0'; ff6c6475433641737731515947564b576b796a6c6b4c773d3d <= (others => '0'); ff566578526b744538644b49392b59753658356a6359413d3d <= ff566578526b744538644b49392b59753658356a6359413d3d + '1'; if (ff566578526b744538644b49392b59753658356a6359413d3d = 255) then if (ff6e3536516f646f71694a6d4152536d735a78574475773d3d /= 0 and ff6e3536516f646f71694a6d4152536d735a78574475773d3d - '1' /= ff6f6f49524b56444d77713077545a545663315a5045413d3d) then ff6f6f49524b56444d77713077545a545663315a5045413d3d <= ff6f6f49524b56444d77713077545a545663315a5045413d3d + '1'; ff70553469356248674669474e4f396e764b594b7958773d3d <= '1'; ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_idle; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '0'; ff566578526b744538644b49392b59753658356a6359413d3d <= (others => '0'); else ff6f6f49524b56444d77713077545a545663315a5045413d3d <= (others => '0'); ff70553469356248674669474e4f396e764b594b7958773d3d <= '0'; ff3332356d7477754d64456339442f2b5a6c44727579413d3d <= st_idle; ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d <= '0'; ff566578526b744538644b49392b59753658356a6359413d3d <= (others => '0'); end if; end if; when others => null; end case; end if; end process; process(ff5265546f48666357584236504c5951756c496d4859773d3d) is begin if rising_edge(ff5265546f48666357584236504c5951756c496d4859773d3d) then if (ff734375372b7345675871315954415046687a5046356b45354d79796e5a506d70346e7835483537776a52733d(0) = '1') then elsif (ff566578526b744538644b49392b59753658356a6359413d3d > 20) then if (ff6e3536516f646f71694a6d4152536d735a78574475773d3d /= 0) then if (ff6e3536516f646f71694a6d4152536d735a78574475773d3d - '1' = ff6f6f49524b56444d77713077545a545663315a5045413d3d) then ff442f5a372f344d4f50427876662b55446d74477771673d3d <= '1'; end if; else ff442f5a372f344d4f50427876662b55446d74477771673d3d <= '1'; end if; end if; end if; end process; process(ff66634b612f4d46776431426239796e69595a575831413d3d) is begin if rising_edge(ff66634b612f4d46776431426239796e69595a575831413d3d) then if (ff734375372b7345675871315954415046687a5046356b45354d79796e5a506d70346e7835483537776a52733d(1) = '1') then elsif (ff526a78674d6b6743434d707672794536766e71794c513d3d = '1') then ff6947484f5a464e57314e6d57485976714235554f44773d3d <= '1'; end if; end if; end process; ff4f4e713355624a533343352b346e33756246377338673d3d <= ff5a6c666e34314c507a4e595439584b4e644d6f326e773d3d; ff78367278306164782f62776f386552346a615a594c673d3d <= '1' when (ff764d71614b5443474d507a536f41756f6a356a5638773d3d = '1' and ff70553469356248674669474e4f396e764b594b7958773d3d = '0') else '0'; U_fifo_generator_0 : entity work.fifo_generator_0 PORT map ( clk => ff66634b612f4d46776431426239796e69595a575831413d3d , rst => not ff35486432672f59566a33374f395741557145392b47413d3d , din => ff71444670796c6e74686577476451676d39424a302f513d3d , wr_en => ff556c7542746b515351533838686b37614254365847513d3d , rd_en => ff5343306145363166474e5241315a39645a6a6d4879773d3d , dout => ff49596952527246685a316551654f564e6635662f39413d3d , full => open , empty => open ); U_fifo_generator_1 : entity work.fifo_generator_0 PORT map ( clk => ff66634b612f4d46776431426239796e69595a575831413d3d , rst => not ff35486432672f59566a33374f395741557145392b47413d3d , din => ff557746415069796532515158714d554e6632366b38513d3d , wr_en => ff74434b38614a354247676547696a3048776554796f513d3d , rd_en => ff4a644751576c526f685a63496b69594a7172304848673d3d , dout => ff644e52654c42493575715935704d6a745041723146773d3d , full => open , empty => open ); ff714f412b3968364e7561522b464c4e355a4a445231673d3d <= ff6d79702b36614f2b55594a797369344e6c56482b65413d3d when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 0) else ff2f4636662f6c3072673535706e41485a3762646854513d3d(16 downto 5) when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 32) else ff2f4636662f6c3072673535706e41485a3762646854513d3d(15 downto 4) when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 16) else ff2f4636662f6c3072673535706e41485a3762646854513d3d(14 downto 3) when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 8) else ff2f4636662f6c3072673535706e41485a3762646854513d3d(13 downto 2) when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 4) else ff2f4636662f6c3072673535706e41485a3762646854513d3d(12 downto 1) when (ff6e3536516f646f71694a6d4152536d735a78574475773d3d = 2); U_DP_RAM : entity work.DP_RAM PORT map ( clka => ff66634b612f4d46776431426239796e69595a575831413d3d, wea => ff366e677746596c337243586a4d5452644a775a4c65673d3d, addra => ff6c6475433641737731515947564b576b796a6c6b4c773d3d, dina => "0000" & ff714f412b3968364e7561522b464c4e355a4a445231673d3d, douta => open, clkb => ff5265546f48666357584236504c5951756c496d4859773d3d, web => "0", addrb => ff41734f64796e456c5746356d69726979457351574d513d3d, dinb => (others=>'0'), doutb => ff71696d73453179677739397a633754775874385361773d3d ); process(ff5265546f48666357584236504c5951756c496d4859773d3d) is begin if rising_edge(ff5265546f48666357584236504c5951756c496d4859773d3d) then ff545336484f3169516e614c77456c316d622f53482f673d3d <= ff35345579546249415444475676365976357270794f706466634b6948397a6f7466675938636851536461593d; if (ff734375372b7345675871315954415046687a5046356b45354d79796e5a506d70346e7835483537776a52733d(0) = '1') then ff41734f64796e456c5746356d69726979457351574d513d3d <= (others=>'0'); ff64684b35757841614e684d304243786e335a6a5438513d3d <= (others => '0'); elsif (ff35345579546249415444475676365976357270794f706466634b6948397a6f7466675938636851536461593d = '1' and ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d = '0') then ff41734f64796e456c5746356d69726979457351574d513d3d <= ff41734f64796e456c5746356d69726979457351574d513d3d + '1'; if (ff507a534d467a36562f345a534e5755745574326668773d3d(0) = '0') then ff64684b35757841614e684d304243786e335a6a5438513d3d(11 downto 0) <= ff64684b35757841614e684d304243786e335a6a5438513d3d(11 downto 0) + '1'; else ff64684b35757841614e684d304243786e335a6a5438513d3d <= ff71696d73453179677739397a633754775874385361773d3d; end if; elsif (ff35345579546249415444475676365976357270794f754e5335735975446a484354684b506d6d344f6554453d = '1' and ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d = '0') then ff41734f64796e456c5746356d69726979457351574d513d3d <= ff41734f64796e456c5746356d69726979457351574d513d3d - '1'; ff64684b35757841614e684d304243786e335a6a5438513d3d(11 downto 0) <= ff64684b35757841614e684d304243786e335a6a5438513d3d(11 downto 0) - '1'; end if; end if; end process; process(ff5265546f48666357584236504c5951756c496d4859773d3d) is begin if rising_edge(ff5265546f48666357584236504c5951756c496d4859773d3d) then if (ff734375372b7345675871315954415046687a5046356b45354d79796e5a506d70346e7835483537776a52733d(1) = '1') then ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d <= x"FFFF"; elsif (ff35345579546249415444475676365976357270794f706466634b6948397a6f7466675938636851536461593d = '1' and ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d = '1') then ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d(11 downto 0) <= ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d(11 downto 0) - '1'; elsif (ff35345579546249415444475676365976357270794f754e5335735975446a484354684b506d6d344f6554453d = '1' and ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d = '1') then ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d(11 downto 0) <= ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d(11 downto 0) + '1'; end if; end if; end process; ff336c46794e7a665a41773233795930316930313174513d3d <= ff537a6f52416d624a366b395532676b7071435155555a6466634b6948397a6f7466675938636851536461593d when (ff4732345242474976646c354951705765616f3543544b68324e585352362b4c533254566936366b482f516f3d = '1') else ff64684b35757841614e684d304243786e335a6a5438513d3d; ff547151597569774e3243584579796a57764a7a6c39673d3d <= ff442f5a372f344d4f50427876662b55446d74477771673d3d; ff3749554e2f736346657730416b38716a732b745371513d3d <= ff6947484f5a464e57314e6d57485976714235554f44773d3d; end Behavioral;