library IEEE; use IEEE.STD_LOGIC_1164.ALL; use IEEE.STD_LOGIC_arith.ALL; use IEEE.STD_LOGIC_unsigned.ALL; library UNISIM; use UNISIM.VComponents.all; use work.pkg_util.all; entity QuadDemod is Port ( ff5178416e525134735a5578472f567a565a2b677774513d3d : in std_logic; ff726531644c73452f3079714267764a6a697277334d413d3d : in std_logic_vector(13 downto 0); ff574a4976744f65433044753745544c46716d417944413d3d : in std_logic_vector(21 downto 0); ff6c6a5873626b4c7468497a6d50736777574234572b673d3d : out std_logic; ff3173395850624f7175547232346b397971375a6f37413d3d : out std_logic_vector(15 downto 0); ff69564244526f7a527376554b6668394a4b6f336b32513d3d : out std_logic_vector(15 downto 0) ); end QuadDemod; architecture Behavioral of QuadDemod is component sincos is Port ( ff5178416e525134735a5578472f567a565a2b677774513d3d : in std_logic; m_reset : in std_logic; m_ce : in std_logic; m_step : in std_logic_vector(21 downto 0); m_cos : out std_logic_vector(15 downto 0); m_sin : out std_logic_vector(15 downto 0)); end component; component sincosNew is Port ( ff5178416e525134735a5578472f567a565a2b677774513d3d : in std_logic; m_step : in std_logic_vector(21 downto 0); m_cos : out std_logic_vector(15 downto 0); m_sin : out std_logic_vector(15 downto 0)); end component; COMPONENT ip_mult_s14_s16 PORT ( CLK : IN STD_LOGIC; A : IN STD_LOGIC_VECTOR(13 DOWNTO 0); B : IN STD_LOGIC_VECTOR(15 DOWNTO 0); P : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) ); END COMPONENT; COMPONENT ip_fifo_adc_din PORT ( wr_clk : IN STD_LOGIC; rd_clk : IN STD_LOGIC; din : IN STD_LOGIC_VECTOR(13 DOWNTO 0); wr_en : IN STD_LOGIC; rd_en : IN STD_LOGIC; dout : OUT STD_LOGIC_VECTOR(13 DOWNTO 0); full : OUT STD_LOGIC; empty : OUT STD_LOGIC ); END COMPONENT; COMPONENT ip_quad_lpf PORT ( aclk : IN STD_LOGIC; s_axis_data_tvalid : IN STD_LOGIC; s_axis_data_tready : OUT STD_LOGIC; s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0); m_axis_data_tvalid : OUT STD_LOGIC; m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0) ); END COMPONENT; signal ff3136724c6d546f35755954616e5959735776315034673d3d : std_logic_vector(13 downto 0); signal ff6664536151446532395630594b7176672f31463342673d3d : std_logic_vector(15 downto 0); signal ff653177574354633548714b463064433133334e4b6c513d3d : std_logic_vector(15 downto 0); signal ff636f2b495a3144664465442b722b4d4a5a4e596857773d3d : std_logic_vector(15 downto 0); signal ff6a7a434e716c7a746f717743306b6f714e6d447a73673d3d : std_logic_vector(15 downto 0); signal ff3938384f57416d52426b7367535242306b696e7962773d3d : std_logic_vector(15 downto 0); signal ff2b4f33497435594648796245634a48454378704c53413d3d : STD_LOGIC_VECTOR(31 DOWNTO 0); signal ff566f39426c6f54753770733169365356423742684e773d3d : STD_LOGIC; signal ff487833466a537a722f5a6d34447563522f4e4e7538413d3d : STD_LOGIC_VECTOR(47 DOWNTO 0); signal ff68695269376a776552687a703771676e4b7a564768773d3d : std_logic_vector(21 downto 0); signal ff767641446948317936577661646545395a44673268513d3d : std_logic; signal ff347675484466586c4e5134582f55506b7837723237413d3d : STD_LOGIC; signal ff4268717a775148596e716545416569594745686f64413d3d : std_logic_vector(15 downto 0); signal ff736f384947544c6f6c545356674e54614361726e69673d3d : std_logic_vector(15 downto 0); COMPONENT ila_qmod PORT ( clk : IN STD_LOGIC; probe0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); probe1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); probe2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); probe3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0)); END COMPONENT ; signal ff6e582f56416e6b615837436b76752f5a756a79724a673d3d : std_logic_vector(15 downto 0); signal ff75417537664168364c76687674384d494559684974513d3d : std_logic_vector(15 downto 0); signal ff6e35716d4d333743366a317539723277426a544356513d3d : std_logic_vector(15 downto 0); signal ff786239515958776d716b30317a70482f516456536c673d3d : std_logic_vector(15 downto 0); begin U_sincosNew : sincosNew Port map( ff5178416e525134735a5578472f567a565a2b677774513d3d => ff5178416e525134735a5578472f567a565a2b677774513d3d , m_step => ff574a4976744f65433044753745544c46716d417944413d3d , m_cos => ff653177574354633548714b463064433133334e4b6c513d3d , m_sin => ff6664536151446532395630594b7176672f31463342673d3d ); inst_i_mult : ip_mult_s14_s16 PORT map( CLK => ff5178416e525134735a5578472f567a565a2b677774513d3d, A => ff726531644c73452f3079714267764a6a697277334d413d3d, B => ff6664536151446532395630594b7176672f31463342673d3d, P => ff6a7a434e716c7a746f717743306b6f714e6d447a73673d3d ); inst_q_mult : ip_mult_s14_s16 PORT map( CLK => ff5178416e525134735a5578472f567a565a2b677774513d3d, A => ff726531644c73452f3079714267764a6a697277334d413d3d, B => ff636f2b495a3144664465442b722b4d4a5a4e596857773d3d, P => ff3938384f57416d52426b7367535242306b696e7962773d3d ); ff636f2b495a3144664465442b722b4d4a5a4e596857773d3d <= not(ff653177574354633548714b463064433133334e4b6c513d3d) + '1'; inst_ip_quad_lpf : ip_quad_lpf PORT map( aclk => ff5178416e525134735a5578472f567a565a2b677774513d3d, s_axis_data_tvalid => '1', s_axis_data_tready => ff767641446948317936577661646545395a44673268513d3d, s_axis_data_tdata => ff2b4f33497435594648796245634a48454378704c53413d3d, m_axis_data_tvalid => ff566f39426c6f54753770733169365356423742684e773d3d, m_axis_data_tdata => ff487833466a537a722f5a6d34447563522f4e4e7538413d3d ); ff2b4f33497435594648796245634a48454378704c53413d3d <= ff6a7a434e716c7a746f717743306b6f714e6d447a73673d3d & ff3938384f57416d52426b7367535242306b696e7962773d3d; process(ff5178416e525134735a5578472f567a565a2b677774513d3d) begin if rising_edge(ff5178416e525134735a5578472f567a565a2b677774513d3d) then ff347675484466586c4e5134582f55506b7837723237413d3d <= ff566f39426c6f54753770733169365356423742684e773d3d; ff4268717a775148596e716545416569594745686f64413d3d <= sat(rnd(ff487833466a537a722f5a6d34447563522f4e4e7538413d3d(47 downto 24),5),3); ff736f384947544c6f6c545356674e54614361726e69673d3d <= sat(rnd(ff487833466a537a722f5a6d34447563522f4e4e7538413d3d(23 downto 0),5),3); end if; end process; process(ff5178416e525134735a5578472f567a565a2b677774513d3d) begin if rising_edge(ff5178416e525134735a5578472f567a565a2b677774513d3d) then ff6c6a5873626b4c7468497a6d50736777574234572b673d3d <= ff347675484466586c4e5134582f55506b7837723237413d3d ; ff3173395850624f7175547232346b397971375a6f37413d3d <= ff4268717a775148596e716545416569594745686f64413d3d ; ff69564244526f7a527376554b6668394a4b6f336b32513d3d <= ff736f384947544c6f6c545356674e54614361726e69673d3d ; end if; end process; end Behavioral;